magic
tech sky130A
magscale 1 2
timestamp 1649709025
<< nwell >>
rect -2915 -864 2915 864
<< pmos >>
rect -2719 -645 -2319 645
rect -2261 -645 -1861 645
rect -1803 -645 -1403 645
rect -1345 -645 -945 645
rect -887 -645 -487 645
rect -429 -645 -29 645
rect 29 -645 429 645
rect 487 -645 887 645
rect 945 -645 1345 645
rect 1403 -645 1803 645
rect 1861 -645 2261 645
rect 2319 -645 2719 645
<< pdiff >>
rect -2777 633 -2719 645
rect -2777 -633 -2765 633
rect -2731 -633 -2719 633
rect -2777 -645 -2719 -633
rect -2319 633 -2261 645
rect -2319 -633 -2307 633
rect -2273 -633 -2261 633
rect -2319 -645 -2261 -633
rect -1861 633 -1803 645
rect -1861 -633 -1849 633
rect -1815 -633 -1803 633
rect -1861 -645 -1803 -633
rect -1403 633 -1345 645
rect -1403 -633 -1391 633
rect -1357 -633 -1345 633
rect -1403 -645 -1345 -633
rect -945 633 -887 645
rect -945 -633 -933 633
rect -899 -633 -887 633
rect -945 -645 -887 -633
rect -487 633 -429 645
rect -487 -633 -475 633
rect -441 -633 -429 633
rect -487 -645 -429 -633
rect -29 633 29 645
rect -29 -633 -17 633
rect 17 -633 29 633
rect -29 -645 29 -633
rect 429 633 487 645
rect 429 -633 441 633
rect 475 -633 487 633
rect 429 -645 487 -633
rect 887 633 945 645
rect 887 -633 899 633
rect 933 -633 945 633
rect 887 -645 945 -633
rect 1345 633 1403 645
rect 1345 -633 1357 633
rect 1391 -633 1403 633
rect 1345 -645 1403 -633
rect 1803 633 1861 645
rect 1803 -633 1815 633
rect 1849 -633 1861 633
rect 1803 -645 1861 -633
rect 2261 633 2319 645
rect 2261 -633 2273 633
rect 2307 -633 2319 633
rect 2261 -645 2319 -633
rect 2719 633 2777 645
rect 2719 -633 2731 633
rect 2765 -633 2777 633
rect 2719 -645 2777 -633
<< pdiffc >>
rect -2765 -633 -2731 633
rect -2307 -633 -2273 633
rect -1849 -633 -1815 633
rect -1391 -633 -1357 633
rect -933 -633 -899 633
rect -475 -633 -441 633
rect -17 -633 17 633
rect 441 -633 475 633
rect 899 -633 933 633
rect 1357 -633 1391 633
rect 1815 -633 1849 633
rect 2273 -633 2307 633
rect 2731 -633 2765 633
<< nsubdiff >>
rect -2879 794 -2783 828
rect 2783 794 2879 828
rect -2879 732 -2845 794
rect 2845 732 2879 794
rect -2879 -794 -2845 -732
rect 2845 -794 2879 -732
rect -2879 -828 -2783 -794
rect 2783 -828 2879 -794
<< nsubdiffcont >>
rect -2783 794 2783 828
rect -2879 -732 -2845 732
rect 2845 -732 2879 732
rect -2783 -828 2783 -794
<< poly >>
rect -2719 726 -2319 742
rect -2719 692 -2703 726
rect -2335 692 -2319 726
rect -2719 645 -2319 692
rect -2261 726 -1861 742
rect -2261 692 -2245 726
rect -1877 692 -1861 726
rect -2261 645 -1861 692
rect -1803 726 -1403 742
rect -1803 692 -1787 726
rect -1419 692 -1403 726
rect -1803 645 -1403 692
rect -1345 726 -945 742
rect -1345 692 -1329 726
rect -961 692 -945 726
rect -1345 645 -945 692
rect -887 726 -487 742
rect -887 692 -871 726
rect -503 692 -487 726
rect -887 645 -487 692
rect -429 726 -29 742
rect -429 692 -413 726
rect -45 692 -29 726
rect -429 645 -29 692
rect 29 726 429 742
rect 29 692 45 726
rect 413 692 429 726
rect 29 645 429 692
rect 487 726 887 742
rect 487 692 503 726
rect 871 692 887 726
rect 487 645 887 692
rect 945 726 1345 742
rect 945 692 961 726
rect 1329 692 1345 726
rect 945 645 1345 692
rect 1403 726 1803 742
rect 1403 692 1419 726
rect 1787 692 1803 726
rect 1403 645 1803 692
rect 1861 726 2261 742
rect 1861 692 1877 726
rect 2245 692 2261 726
rect 1861 645 2261 692
rect 2319 726 2719 742
rect 2319 692 2335 726
rect 2703 692 2719 726
rect 2319 645 2719 692
rect -2719 -692 -2319 -645
rect -2719 -726 -2703 -692
rect -2335 -726 -2319 -692
rect -2719 -742 -2319 -726
rect -2261 -692 -1861 -645
rect -2261 -726 -2245 -692
rect -1877 -726 -1861 -692
rect -2261 -742 -1861 -726
rect -1803 -692 -1403 -645
rect -1803 -726 -1787 -692
rect -1419 -726 -1403 -692
rect -1803 -742 -1403 -726
rect -1345 -692 -945 -645
rect -1345 -726 -1329 -692
rect -961 -726 -945 -692
rect -1345 -742 -945 -726
rect -887 -692 -487 -645
rect -887 -726 -871 -692
rect -503 -726 -487 -692
rect -887 -742 -487 -726
rect -429 -692 -29 -645
rect -429 -726 -413 -692
rect -45 -726 -29 -692
rect -429 -742 -29 -726
rect 29 -692 429 -645
rect 29 -726 45 -692
rect 413 -726 429 -692
rect 29 -742 429 -726
rect 487 -692 887 -645
rect 487 -726 503 -692
rect 871 -726 887 -692
rect 487 -742 887 -726
rect 945 -692 1345 -645
rect 945 -726 961 -692
rect 1329 -726 1345 -692
rect 945 -742 1345 -726
rect 1403 -692 1803 -645
rect 1403 -726 1419 -692
rect 1787 -726 1803 -692
rect 1403 -742 1803 -726
rect 1861 -692 2261 -645
rect 1861 -726 1877 -692
rect 2245 -726 2261 -692
rect 1861 -742 2261 -726
rect 2319 -692 2719 -645
rect 2319 -726 2335 -692
rect 2703 -726 2719 -692
rect 2319 -742 2719 -726
<< polycont >>
rect -2703 692 -2335 726
rect -2245 692 -1877 726
rect -1787 692 -1419 726
rect -1329 692 -961 726
rect -871 692 -503 726
rect -413 692 -45 726
rect 45 692 413 726
rect 503 692 871 726
rect 961 692 1329 726
rect 1419 692 1787 726
rect 1877 692 2245 726
rect 2335 692 2703 726
rect -2703 -726 -2335 -692
rect -2245 -726 -1877 -692
rect -1787 -726 -1419 -692
rect -1329 -726 -961 -692
rect -871 -726 -503 -692
rect -413 -726 -45 -692
rect 45 -726 413 -692
rect 503 -726 871 -692
rect 961 -726 1329 -692
rect 1419 -726 1787 -692
rect 1877 -726 2245 -692
rect 2335 -726 2703 -692
<< locali >>
rect -2879 794 -2783 828
rect 2783 794 2879 828
rect -2879 732 -2845 794
rect 2845 732 2879 794
rect -2719 692 -2703 726
rect -2335 692 -2319 726
rect -2261 692 -2245 726
rect -1877 692 -1861 726
rect -1803 692 -1787 726
rect -1419 692 -1403 726
rect -1345 692 -1329 726
rect -961 692 -945 726
rect -887 692 -871 726
rect -503 692 -487 726
rect -429 692 -413 726
rect -45 692 -29 726
rect 29 692 45 726
rect 413 692 429 726
rect 487 692 503 726
rect 871 692 887 726
rect 945 692 961 726
rect 1329 692 1345 726
rect 1403 692 1419 726
rect 1787 692 1803 726
rect 1861 692 1877 726
rect 2245 692 2261 726
rect 2319 692 2335 726
rect 2703 692 2719 726
rect -2765 633 -2731 649
rect -2765 -649 -2731 -633
rect -2307 633 -2273 649
rect -2307 -649 -2273 -633
rect -1849 633 -1815 649
rect -1849 -649 -1815 -633
rect -1391 633 -1357 649
rect -1391 -649 -1357 -633
rect -933 633 -899 649
rect -933 -649 -899 -633
rect -475 633 -441 649
rect -475 -649 -441 -633
rect -17 633 17 649
rect -17 -649 17 -633
rect 441 633 475 649
rect 441 -649 475 -633
rect 899 633 933 649
rect 899 -649 933 -633
rect 1357 633 1391 649
rect 1357 -649 1391 -633
rect 1815 633 1849 649
rect 1815 -649 1849 -633
rect 2273 633 2307 649
rect 2273 -649 2307 -633
rect 2731 633 2765 649
rect 2731 -649 2765 -633
rect -2719 -726 -2703 -692
rect -2335 -726 -2319 -692
rect -2261 -726 -2245 -692
rect -1877 -726 -1861 -692
rect -1803 -726 -1787 -692
rect -1419 -726 -1403 -692
rect -1345 -726 -1329 -692
rect -961 -726 -945 -692
rect -887 -726 -871 -692
rect -503 -726 -487 -692
rect -429 -726 -413 -692
rect -45 -726 -29 -692
rect 29 -726 45 -692
rect 413 -726 429 -692
rect 487 -726 503 -692
rect 871 -726 887 -692
rect 945 -726 961 -692
rect 1329 -726 1345 -692
rect 1403 -726 1419 -692
rect 1787 -726 1803 -692
rect 1861 -726 1877 -692
rect 2245 -726 2261 -692
rect 2319 -726 2335 -692
rect 2703 -726 2719 -692
rect -2879 -794 -2845 -732
rect 2845 -794 2879 -732
rect -2879 -828 -2783 -794
rect 2783 -828 2879 -794
<< viali >>
rect -2703 692 -2335 726
rect -2245 692 -1877 726
rect -1787 692 -1419 726
rect -1329 692 -961 726
rect -871 692 -503 726
rect -413 692 -45 726
rect 45 692 413 726
rect 503 692 871 726
rect 961 692 1329 726
rect 1419 692 1787 726
rect 1877 692 2245 726
rect 2335 692 2703 726
rect -2765 -633 -2731 633
rect -2307 -633 -2273 633
rect -1849 -633 -1815 633
rect -1391 -633 -1357 633
rect -933 -633 -899 633
rect -475 -633 -441 633
rect -17 -633 17 633
rect 441 -633 475 633
rect 899 -633 933 633
rect 1357 -633 1391 633
rect 1815 -633 1849 633
rect 2273 -633 2307 633
rect 2731 -633 2765 633
rect -2703 -726 -2335 -692
rect -2245 -726 -1877 -692
rect -1787 -726 -1419 -692
rect -1329 -726 -961 -692
rect -871 -726 -503 -692
rect -413 -726 -45 -692
rect 45 -726 413 -692
rect 503 -726 871 -692
rect 961 -726 1329 -692
rect 1419 -726 1787 -692
rect 1877 -726 2245 -692
rect 2335 -726 2703 -692
<< metal1 >>
rect -2715 726 -2323 732
rect -2715 692 -2703 726
rect -2335 692 -2323 726
rect -2715 686 -2323 692
rect -2257 726 -1865 732
rect -2257 692 -2245 726
rect -1877 692 -1865 726
rect -2257 686 -1865 692
rect -1799 726 -1407 732
rect -1799 692 -1787 726
rect -1419 692 -1407 726
rect -1799 686 -1407 692
rect -1341 726 -949 732
rect -1341 692 -1329 726
rect -961 692 -949 726
rect -1341 686 -949 692
rect -883 726 -491 732
rect -883 692 -871 726
rect -503 692 -491 726
rect -883 686 -491 692
rect -425 726 -33 732
rect -425 692 -413 726
rect -45 692 -33 726
rect -425 686 -33 692
rect 33 726 425 732
rect 33 692 45 726
rect 413 692 425 726
rect 33 686 425 692
rect 491 726 883 732
rect 491 692 503 726
rect 871 692 883 726
rect 491 686 883 692
rect 949 726 1341 732
rect 949 692 961 726
rect 1329 692 1341 726
rect 949 686 1341 692
rect 1407 726 1799 732
rect 1407 692 1419 726
rect 1787 692 1799 726
rect 1407 686 1799 692
rect 1865 726 2257 732
rect 1865 692 1877 726
rect 2245 692 2257 726
rect 1865 686 2257 692
rect 2323 726 2715 732
rect 2323 692 2335 726
rect 2703 692 2715 726
rect 2323 686 2715 692
rect -2771 633 -2725 645
rect -2771 -633 -2765 633
rect -2731 -633 -2725 633
rect -2771 -645 -2725 -633
rect -2313 633 -2267 645
rect -2313 -633 -2307 633
rect -2273 -633 -2267 633
rect -2313 -645 -2267 -633
rect -1855 633 -1809 645
rect -1855 -633 -1849 633
rect -1815 -633 -1809 633
rect -1855 -645 -1809 -633
rect -1397 633 -1351 645
rect -1397 -633 -1391 633
rect -1357 -633 -1351 633
rect -1397 -645 -1351 -633
rect -939 633 -893 645
rect -939 -633 -933 633
rect -899 -633 -893 633
rect -939 -645 -893 -633
rect -481 633 -435 645
rect -481 -633 -475 633
rect -441 -633 -435 633
rect -481 -645 -435 -633
rect -23 633 23 645
rect -23 -633 -17 633
rect 17 -633 23 633
rect -23 -645 23 -633
rect 435 633 481 645
rect 435 -633 441 633
rect 475 -633 481 633
rect 435 -645 481 -633
rect 893 633 939 645
rect 893 -633 899 633
rect 933 -633 939 633
rect 893 -645 939 -633
rect 1351 633 1397 645
rect 1351 -633 1357 633
rect 1391 -633 1397 633
rect 1351 -645 1397 -633
rect 1809 633 1855 645
rect 1809 -633 1815 633
rect 1849 -633 1855 633
rect 1809 -645 1855 -633
rect 2267 633 2313 645
rect 2267 -633 2273 633
rect 2307 -633 2313 633
rect 2267 -645 2313 -633
rect 2725 633 2771 645
rect 2725 -633 2731 633
rect 2765 -633 2771 633
rect 2725 -645 2771 -633
rect -2715 -692 -2323 -686
rect -2715 -726 -2703 -692
rect -2335 -726 -2323 -692
rect -2715 -732 -2323 -726
rect -2257 -692 -1865 -686
rect -2257 -726 -2245 -692
rect -1877 -726 -1865 -692
rect -2257 -732 -1865 -726
rect -1799 -692 -1407 -686
rect -1799 -726 -1787 -692
rect -1419 -726 -1407 -692
rect -1799 -732 -1407 -726
rect -1341 -692 -949 -686
rect -1341 -726 -1329 -692
rect -961 -726 -949 -692
rect -1341 -732 -949 -726
rect -883 -692 -491 -686
rect -883 -726 -871 -692
rect -503 -726 -491 -692
rect -883 -732 -491 -726
rect -425 -692 -33 -686
rect -425 -726 -413 -692
rect -45 -726 -33 -692
rect -425 -732 -33 -726
rect 33 -692 425 -686
rect 33 -726 45 -692
rect 413 -726 425 -692
rect 33 -732 425 -726
rect 491 -692 883 -686
rect 491 -726 503 -692
rect 871 -726 883 -692
rect 491 -732 883 -726
rect 949 -692 1341 -686
rect 949 -726 961 -692
rect 1329 -726 1341 -692
rect 949 -732 1341 -726
rect 1407 -692 1799 -686
rect 1407 -726 1419 -692
rect 1787 -726 1799 -692
rect 1407 -732 1799 -726
rect 1865 -692 2257 -686
rect 1865 -726 1877 -692
rect 2245 -726 2257 -692
rect 1865 -732 2257 -726
rect 2323 -692 2715 -686
rect 2323 -726 2335 -692
rect 2703 -726 2715 -692
rect 2323 -732 2715 -726
<< properties >>
string FIXED_BBOX -2862 -811 2862 811
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.45 l 2 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
