magic
tech sky130A
magscale 1 2
timestamp 1649715113
<< nwell >>
rect -2813 -707 2813 707
<< pmos >>
rect -2719 -645 -2319 645
rect -2261 -645 -1861 645
rect -1803 -645 -1403 645
rect -1345 -645 -945 645
rect -887 -645 -487 645
rect -429 -645 -29 645
rect 29 -645 429 645
rect 487 -645 887 645
rect 945 -645 1345 645
rect 1403 -645 1803 645
rect 1861 -645 2261 645
rect 2319 -645 2719 645
<< pdiff >>
rect -2777 633 -2719 645
rect -2777 -633 -2765 633
rect -2731 -633 -2719 633
rect -2777 -645 -2719 -633
rect -2319 633 -2261 645
rect -2319 -633 -2307 633
rect -2273 -633 -2261 633
rect -2319 -645 -2261 -633
rect -1861 633 -1803 645
rect -1861 -633 -1849 633
rect -1815 -633 -1803 633
rect -1861 -645 -1803 -633
rect -1403 633 -1345 645
rect -1403 -633 -1391 633
rect -1357 -633 -1345 633
rect -1403 -645 -1345 -633
rect -945 633 -887 645
rect -945 -633 -933 633
rect -899 -633 -887 633
rect -945 -645 -887 -633
rect -487 633 -429 645
rect -487 -633 -475 633
rect -441 -633 -429 633
rect -487 -645 -429 -633
rect -29 633 29 645
rect -29 -633 -17 633
rect 17 -633 29 633
rect -29 -645 29 -633
rect 429 633 487 645
rect 429 -633 441 633
rect 475 -633 487 633
rect 429 -645 487 -633
rect 887 633 945 645
rect 887 -633 899 633
rect 933 -633 945 633
rect 887 -645 945 -633
rect 1345 633 1403 645
rect 1345 -633 1357 633
rect 1391 -633 1403 633
rect 1345 -645 1403 -633
rect 1803 633 1861 645
rect 1803 -633 1815 633
rect 1849 -633 1861 633
rect 1803 -645 1861 -633
rect 2261 633 2319 645
rect 2261 -633 2273 633
rect 2307 -633 2319 633
rect 2261 -645 2319 -633
rect 2719 633 2777 645
rect 2719 -633 2731 633
rect 2765 -633 2777 633
rect 2719 -645 2777 -633
<< pdiffc >>
rect -2765 -633 -2731 633
rect -2307 -633 -2273 633
rect -1849 -633 -1815 633
rect -1391 -633 -1357 633
rect -933 -633 -899 633
rect -475 -633 -441 633
rect -17 -633 17 633
rect 441 -633 475 633
rect 899 -633 933 633
rect 1357 -633 1391 633
rect 1815 -633 1849 633
rect 2273 -633 2307 633
rect 2731 -633 2765 633
<< poly >>
rect -2719 645 -2319 671
rect -2261 645 -1861 671
rect -1803 645 -1403 671
rect -1345 645 -945 671
rect -887 645 -487 671
rect -429 645 -29 671
rect 29 645 429 671
rect 487 645 887 671
rect 945 645 1345 671
rect 1403 645 1803 671
rect 1861 645 2261 671
rect 2319 645 2719 671
rect -2719 -671 -2319 -645
rect -2261 -671 -1861 -645
rect -1803 -671 -1403 -645
rect -1345 -671 -945 -645
rect -887 -671 -487 -645
rect -429 -671 -29 -645
rect 29 -671 429 -645
rect 487 -671 887 -645
rect 945 -671 1345 -645
rect 1403 -671 1803 -645
rect 1861 -671 2261 -645
rect 2319 -671 2719 -645
<< locali >>
rect -2765 633 -2731 649
rect -2765 -649 -2731 -633
rect -2307 633 -2273 649
rect -2307 -649 -2273 -633
rect -1849 633 -1815 649
rect -1849 -649 -1815 -633
rect -1391 633 -1357 649
rect -1391 -649 -1357 -633
rect -933 633 -899 649
rect -933 -649 -899 -633
rect -475 633 -441 649
rect -475 -649 -441 -633
rect -17 633 17 649
rect -17 -649 17 -633
rect 441 633 475 649
rect 441 -649 475 -633
rect 899 633 933 649
rect 899 -649 933 -633
rect 1357 633 1391 649
rect 1357 -649 1391 -633
rect 1815 633 1849 649
rect 1815 -649 1849 -633
rect 2273 633 2307 649
rect 2273 -649 2307 -633
rect 2731 633 2765 649
rect 2731 -649 2765 -633
<< viali >>
rect -2765 -506 -2731 506
rect -2307 -506 -2273 506
rect -1849 -506 -1815 506
rect -1391 -506 -1357 506
rect -933 -506 -899 506
rect -475 -506 -441 506
rect -17 -506 17 506
rect 441 -506 475 506
rect 899 -506 933 506
rect 1357 -506 1391 506
rect 1815 -506 1849 506
rect 2273 -506 2307 506
rect 2731 -506 2765 506
<< metal1 >>
rect -2771 506 -2725 518
rect -2771 -506 -2765 506
rect -2731 -506 -2725 506
rect -2771 -518 -2725 -506
rect -2313 506 -2267 518
rect -2313 -506 -2307 506
rect -2273 -506 -2267 506
rect -2313 -518 -2267 -506
rect -1855 506 -1809 518
rect -1855 -506 -1849 506
rect -1815 -506 -1809 506
rect -1855 -518 -1809 -506
rect -1397 506 -1351 518
rect -1397 -506 -1391 506
rect -1357 -506 -1351 506
rect -1397 -518 -1351 -506
rect -939 506 -893 518
rect -939 -506 -933 506
rect -899 -506 -893 506
rect -939 -518 -893 -506
rect -481 506 -435 518
rect -481 -506 -475 506
rect -441 -506 -435 506
rect -481 -518 -435 -506
rect -23 506 23 518
rect -23 -506 -17 506
rect 17 -506 23 506
rect -23 -518 23 -506
rect 435 506 481 518
rect 435 -506 441 506
rect 475 -506 481 506
rect 435 -518 481 -506
rect 893 506 939 518
rect 893 -506 899 506
rect 933 -506 939 506
rect 893 -518 939 -506
rect 1351 506 1397 518
rect 1351 -506 1357 506
rect 1391 -506 1397 506
rect 1351 -518 1397 -506
rect 1809 506 1855 518
rect 1809 -506 1815 506
rect 1849 -506 1855 506
rect 1809 -518 1855 -506
rect 2267 506 2313 518
rect 2267 -506 2273 506
rect 2307 -506 2313 506
rect 2267 -518 2313 -506
rect 2725 506 2771 518
rect 2725 -506 2731 506
rect 2765 -506 2771 506
rect 2725 -518 2771 -506
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.45 l 2 m 1 nf 12 diffcov 100 polycov 80 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 0 rlcov 0 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 80 viadrn 80 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
