magic
tech sky130A
magscale 1 2
timestamp 1649753498
<< poly >>
rect -2572 -816 -2452 -646
rect -2116 -816 -1996 -646
rect -1660 -816 -1540 -646
rect -1204 -816 -1084 -646
rect -748 -816 -628 -646
rect -292 -816 -172 -646
rect 164 -816 284 -646
rect 620 -816 740 -646
rect 1076 -816 1196 -646
rect 1532 -816 1652 -646
rect 1988 -816 2108 -646
rect 2444 -816 2564 -646
rect -2812 -836 2812 -816
rect -2812 -896 -2642 -836
rect -2582 -896 -2242 -836
rect -2182 -896 -1842 -836
rect -1782 -896 -1442 -836
rect -1382 -896 -1042 -836
rect -982 -896 -642 -836
rect -582 -896 -242 -836
rect -182 -896 158 -836
rect 218 -896 558 -836
rect 618 -896 958 -836
rect 1018 -896 1358 -836
rect 1418 -896 1758 -836
rect 1818 -896 2158 -836
rect 2218 -896 2558 -836
rect 2618 -896 2812 -836
rect -2812 -916 2812 -896
<< polycont >>
rect -2642 -896 -2582 -836
rect -2242 -896 -2182 -836
rect -1842 -896 -1782 -836
rect -1442 -896 -1382 -836
rect -1042 -896 -982 -836
rect -642 -896 -582 -836
rect -242 -896 -182 -836
rect 158 -896 218 -836
rect 558 -896 618 -836
rect 958 -896 1018 -836
rect 1358 -896 1418 -836
rect 1758 -896 1818 -836
rect 2158 -896 2218 -836
rect 2558 -896 2618 -836
<< locali >>
rect -2812 850 -2642 910
rect -2582 850 -2242 910
rect -2182 850 -1842 910
rect -1782 850 -1442 910
rect -1382 850 -1042 910
rect -982 850 -642 910
rect -582 850 -242 910
rect -182 850 158 910
rect 218 850 558 910
rect 618 850 958 910
rect 1018 850 1358 910
rect 1418 850 1758 910
rect 1818 850 2158 910
rect 2218 850 2558 910
rect 2618 850 2812 910
rect -2812 730 2812 790
rect -2308 626 -2274 730
rect -1392 626 -1358 730
rect -476 626 -442 730
rect 440 626 474 730
rect 1356 626 1390 730
rect 2272 626 2306 730
rect -2766 -730 -2732 -626
rect -1850 -730 -1816 -626
rect -934 -730 -900 -626
rect -18 -730 16 -626
rect 898 -730 932 -626
rect 1814 -730 1848 -626
rect 2730 -730 2764 -626
rect -2812 -790 2812 -730
rect -2812 -896 -2642 -836
rect -2582 -896 -2242 -836
rect -2182 -896 -1842 -836
rect -1782 -896 -1442 -836
rect -1382 -896 -1042 -836
rect -982 -896 -642 -836
rect -582 -896 -242 -836
rect -182 -896 158 -836
rect 218 -896 558 -836
rect 618 -896 958 -836
rect 1018 -896 1358 -836
rect 1418 -896 1758 -836
rect 1818 -896 2158 -836
rect 2218 -896 2558 -836
rect 2618 -896 2812 -836
rect -2812 -1030 -2642 -970
rect -2582 -1030 -2242 -970
rect -2182 -1030 -1842 -970
rect -1782 -1030 -1442 -970
rect -1382 -1030 -1042 -970
rect -982 -1030 -642 -970
rect -582 -1030 -242 -970
rect -182 -1030 158 -970
rect 218 -1030 558 -970
rect 618 -1030 958 -970
rect 1018 -1030 1358 -970
rect 1418 -1030 1758 -970
rect 1818 -1030 2158 -970
rect 2218 -1030 2558 -970
rect 2618 -1030 2812 -970
<< viali >>
rect -2642 850 -2582 910
rect -2242 850 -2182 910
rect -1842 850 -1782 910
rect -1442 850 -1382 910
rect -1042 850 -982 910
rect -642 850 -582 910
rect -242 850 -182 910
rect 158 850 218 910
rect 558 850 618 910
rect 958 850 1018 910
rect 1358 850 1418 910
rect 1758 850 1818 910
rect 2158 850 2218 910
rect 2558 850 2618 910
rect -2642 -1030 -2582 -970
rect -2242 -1030 -2182 -970
rect -1842 -1030 -1782 -970
rect -1442 -1030 -1382 -970
rect -1042 -1030 -982 -970
rect -642 -1030 -582 -970
rect -242 -1030 -182 -970
rect 158 -1030 218 -970
rect 558 -1030 618 -970
rect 958 -1030 1018 -970
rect 1358 -1030 1418 -970
rect 1758 -1030 1818 -970
rect 2158 -1030 2218 -970
rect 2558 -1030 2618 -970
<< metal1 >>
rect -2812 910 2812 940
rect -2812 850 -2642 910
rect -2582 850 -2242 910
rect -2182 850 -1842 910
rect -1782 850 -1442 910
rect -1382 850 -1042 910
rect -982 850 -642 910
rect -582 850 -242 910
rect -182 850 158 910
rect 218 850 558 910
rect 618 850 958 910
rect 1018 850 1358 910
rect 1418 850 1758 910
rect 1818 850 2158 910
rect 2218 850 2558 910
rect 2618 850 2812 910
rect -2812 820 2812 850
rect -2812 -970 2812 -940
rect -2812 -1030 -2642 -970
rect -2582 -1030 -2242 -970
rect -2182 -1030 -1842 -970
rect -1782 -1030 -1442 -970
rect -1382 -1030 -1042 -970
rect -982 -1030 -642 -970
rect -582 -1030 -242 -970
rect -182 -1030 158 -970
rect 218 -1030 558 -970
rect 618 -1030 958 -970
rect 1018 -1030 1358 -970
rect 1418 -1030 1758 -970
rect 1818 -1030 2158 -970
rect 2218 -1030 2558 -970
rect 2618 -1030 2812 -970
rect -2812 -1060 2812 -1030
use sky130_fd_pr__pfet_01v8_lvt_5AFWP4  xm1
timestamp 0
transform 1 0 0 0 1 0
box -2813 -707 2813 707
<< labels >>
flabel metal1 -2812 850 -2752 910 1 FreeSans 480 0 0 0 VDD
flabel metal1 -2812 -1030 -2752 -970 1 FreeSans 480 0 0 0 VSS
flabel locali 2752 730 2812 790 1 FreeSans 480 0 0 0 SOURCE
flabel locali 2752 -790 2812 -730 1 FreeSans 480 0 0 0 DRAIN
flabel locali 2752 -896 2812 -836 1 FreeSans 480 0 0 0 GATE
<< end >>
