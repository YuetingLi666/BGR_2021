magic
tech sky130A
magscale 1 2
timestamp 1649753335
<< poly >>
rect -2570 -536 -2450 -366
rect -2114 -536 -1994 -366
rect -1658 -536 -1538 -366
rect -1202 -536 -1082 -366
rect -746 -536 -626 -366
rect -290 -536 -170 -366
rect 166 -536 286 -366
rect 622 -536 742 -366
rect 1078 -536 1198 -366
rect 1534 -536 1654 -366
rect 1990 -536 2110 -366
rect 2446 -536 2566 -366
rect -2776 -556 2776 -536
rect -2776 -616 -2606 -556
rect -2546 -616 -2206 -556
rect -2146 -616 -1806 -556
rect -1746 -616 -1406 -556
rect -1346 -616 -1006 -556
rect -946 -616 -606 -556
rect -546 -616 -206 -556
rect -146 -616 194 -556
rect 254 -616 594 -556
rect 654 -616 994 -556
rect 1054 -616 1394 -556
rect 1454 -616 1794 -556
rect 1854 -616 2194 -556
rect 2254 -616 2594 -556
rect 2654 -616 2776 -556
rect -2776 -636 2776 -616
<< polycont >>
rect -2606 -616 -2546 -556
rect -2206 -616 -2146 -556
rect -1806 -616 -1746 -556
rect -1406 -616 -1346 -556
rect -1006 -616 -946 -556
rect -606 -616 -546 -556
rect -206 -616 -146 -556
rect 194 -616 254 -556
rect 594 -616 654 -556
rect 994 -616 1054 -556
rect 1394 -616 1454 -556
rect 1794 -616 1854 -556
rect 2194 -616 2254 -556
rect 2594 -616 2654 -556
<< locali >>
rect -2776 850 -2606 910
rect -2546 850 -2206 910
rect -2146 850 -1806 910
rect -1746 850 -1406 910
rect -1346 850 -1006 910
rect -946 850 -606 910
rect -546 850 -206 910
rect -146 850 194 910
rect 254 850 594 910
rect 654 850 994 910
rect 1054 850 1394 910
rect 1454 850 1794 910
rect 1854 850 2194 910
rect 2254 850 2594 910
rect 2654 850 2776 910
rect -2776 730 2776 790
rect -2306 346 -2272 730
rect -1390 346 -1356 730
rect -474 346 -440 730
rect 442 346 476 730
rect 1358 346 1392 730
rect 2274 346 2308 730
rect -2764 -556 -2730 -346
rect -1848 -556 -1814 -346
rect -932 -556 -898 -346
rect -16 -556 18 -346
rect 900 -556 934 -346
rect 1816 -556 1850 -346
rect -2776 -616 -2606 -556
rect -2546 -616 -2206 -556
rect -2146 -616 -1806 -556
rect -1746 -616 -1406 -556
rect -1346 -616 -1006 -556
rect -946 -616 -606 -556
rect -546 -616 -206 -556
rect -146 -616 194 -556
rect 254 -616 594 -556
rect 654 -616 994 -556
rect 1054 -616 1394 -556
rect 1454 -616 1794 -556
rect 1854 -616 2194 -556
rect 2254 -616 2594 -556
rect 2654 -616 2776 -556
rect -2764 -730 -2730 -616
rect -1848 -730 -1814 -616
rect -932 -730 -898 -616
rect -16 -730 18 -616
rect 900 -730 934 -616
rect 1816 -730 1850 -616
rect -2776 -790 2776 -730
rect -2776 -1030 -2606 -970
rect -2546 -1030 -2206 -970
rect -2146 -1030 -1806 -970
rect -1746 -1030 -1406 -970
rect -1346 -1030 -1006 -970
rect -946 -1030 -606 -970
rect -546 -1030 -206 -970
rect -146 -1030 194 -970
rect 254 -1030 594 -970
rect 654 -1030 994 -970
rect 1054 -1030 1394 -970
rect 1454 -1030 1794 -970
rect 1854 -1030 2194 -970
rect 2254 -1030 2594 -970
rect 2654 -1030 2776 -970
<< viali >>
rect -2606 850 -2546 910
rect -2206 850 -2146 910
rect -1806 850 -1746 910
rect -1406 850 -1346 910
rect -1006 850 -946 910
rect -606 850 -546 910
rect -206 850 -146 910
rect 194 850 254 910
rect 594 850 654 910
rect 994 850 1054 910
rect 1394 850 1454 910
rect 1794 850 1854 910
rect 2194 850 2254 910
rect 2594 850 2654 910
rect -2606 -1030 -2546 -970
rect -2206 -1030 -2146 -970
rect -1806 -1030 -1746 -970
rect -1406 -1030 -1346 -970
rect -1006 -1030 -946 -970
rect -606 -1030 -546 -970
rect -206 -1030 -146 -970
rect 194 -1030 254 -970
rect 594 -1030 654 -970
rect 994 -1030 1054 -970
rect 1394 -1030 1454 -970
rect 1794 -1030 1854 -970
rect 2194 -1030 2254 -970
rect 2594 -1030 2654 -970
<< metal1 >>
rect -2776 910 2776 940
rect -2776 850 -2606 910
rect -2546 850 -2206 910
rect -2146 850 -1806 910
rect -1746 850 -1406 910
rect -1346 850 -1006 910
rect -946 850 -606 910
rect -546 850 -206 910
rect -146 850 194 910
rect 254 850 594 910
rect 654 850 994 910
rect 1054 850 1394 910
rect 1454 850 1794 910
rect 1854 850 2194 910
rect 2254 850 2594 910
rect 2654 850 2776 910
rect -2776 820 2776 850
rect -2776 -970 2776 -940
rect -2776 -1030 -2606 -970
rect -2546 -1030 -2206 -970
rect -2146 -1030 -1806 -970
rect -1746 -1030 -1406 -970
rect -1346 -1030 -1006 -970
rect -946 -1030 -606 -970
rect -546 -1030 -206 -970
rect -146 -1030 194 -970
rect 254 -1030 594 -970
rect 654 -1030 994 -970
rect 1054 -1030 1394 -970
rect 1454 -1030 1794 -970
rect 1854 -1030 2194 -970
rect 2254 -1030 2594 -970
rect 2654 -1030 2776 -970
rect -2776 -1060 2776 -1030
use sky130_fd_pr__nfet_01v8_lvt_UH36AP  xm1
timestamp 0
transform 1 0 0 0 1 0
box -2777 -426 2777 426
<< labels >>
flabel metal1 -2776 850 -2716 910 1 FreeSans 480 0 0 0 VDD
flabel metal1 -2776 -1030 -2716 -970 1 FreeSans 480 0 0 0 VSS
flabel locali 2716 730 2776 790 1 FreeSans 480 0 0 0 SOURCE
flabel locali 2716 -790 2776 -730 1 FreeSans 480 0 0 0 DRAIN
flabel locali 2716 -616 2776 -556 1 FreeSans 480 0 0 0 GATE
<< end >>
